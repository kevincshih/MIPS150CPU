module UATransmit(
  input   Clock,
  input   Reset,

  input   [7:0] DataIn,
  input         DataInValid,
  output        DataInReady,

  output        SOut
);
  // for log2 function
  `include "util.vh"

  //--|Parameters|--------------------------------------------------------------

  parameter   ClockFreq         =   100_000_000;
  parameter   BaudRate          =   115_200;

  // See diagram in the lab guide
  localparam  SymbolEdgeTime    =   ClockFreq / BaudRate;
  localparam  ClockCounterWidth =   log2(SymbolEdgeTime);

  //--|Solution|----------------------------------------------------------------

  wire                            SymbolEdge;
  wire                            Start;
  wire                            TXRunning;

  reg     [3:0]                   BitCounter;
  reg     [ClockCounterWidth-1:0] ClockCounter;
  reg 				  Temp;

  assign DataInReady = ~TXRunning;
  assign Start = DataInValid && DataInReady;
  assign  SymbolEdge   = (ClockCounter == SymbolEdgeTime - 1);
  assign TXRunning = ~(BitCounter == 0);
  assign SOut = Temp;

  // Counts cycles until a single symbol is done
  always @ (posedge Clock) begin
    ClockCounter <= (Start || Reset || SymbolEdge) ? 0 : ClockCounter + 1;
  end

  // Counts down from 10 bits for every character
  always @ (posedge Clock) begin
    if (Reset) begin
      BitCounter <= 0;
    end else if (Start) begin
      BitCounter <= 10;
    end else if (SymbolEdge && TXRunning) begin
      BitCounter <= BitCounter - 1;
    end
  end

  always @ (posedge Clock) begin
    if (TXRunning) begin
	if(BitCounter == 10) Temp <= 1'b0;
	else if (BitCounter == 1) Temp <= 1'b1;
	else Temp <= DataIn[9 - BitCounter];
	end
    else Temp = 1'b1;
  end

endmodule
