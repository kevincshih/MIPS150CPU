module	sar(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			TB,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			D,
			EOC
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					TB;
	//input enter;
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output	   [9:0] D;
	output				EOC;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	localparam
	      S_0 = 4'd0,
		    S_1 = 4'd1,
		    S_2 = 4'd2,
		    S_3 = 4'd3,
		    S_4 = 4'd4,
		    S_5 = 4'd5,
		    S_6 = 4'd6,
		    S_7 = 4'd7,
		    S_8 = 4'd8,
		    Done = 4'd9;
		    
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	wire tb;
	//reg [9:0] out;
	reg d0, d1, d2, d3, d4, d5, d6, d7, d8, d9;
	reg [3:0] CurrentState;
	reg [3:0] NextState;

	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------
	assign tb = TB;
	assign D = {d0, d1, d2, d3, d4, d5, d6, d7, d8, d9};
	assign EOC = (CurrentState == Done);
	
	always@(posedge Clock) begin
	  if (Reset) begin
	     CurrentState <= S_0;
	     {d0,d1,d2,d3,d4,d5,d6,d7,d8,d9} <= 10'd0;
	     //out <= 10'd0;
	     end
	  else CurrentState <= NextState;
	end

	always@(*) begin
		NextState = CurrentState;
		if (Clock) begin
		case(NextState)
		    S_0: begin 
		      d0 = (TB) ? 0 : 1;
		      NextState = S_1;
		      end
		    S_1: begin 
		      d1 = (TB) ? 0 : 1;
		      NextState = S_2;
		      end
		    S_2: begin 
		      d2 = (TB) ? 0 : 1;
		      NextState = S_3;
		      end
		    S_3: begin 
		      d3 = (TB) ? 0 : 1;
		      NextState = S_4;
		      end
		    S_4: begin 
		      d4 = (TB) ? 0 : 1;
		      NextState = S_5;
		      end
		    S_5: begin 
		      d5 = (TB) ? 0 : 1;
		      NextState = S_6;
		      end
		    S_6: begin 
		      d6 = (TB) ? 0 : 1;
		      NextState = S_7;
		      end
		    S_7: begin 
		      d7 = (TB) ? 0 : 1;
		      NextState = S_8;
		      end
		    S_8: begin 
		      d8 = (TB) ? 0 : 1;
		      NextState = Done;
		      end
		    Done: begin 
		      d9 = (TB) ? 0 : 1;
		      //out = {d0,d1,d2,d3,d4,d5,d6,d7,d8,d9}
		      NextState = Done;
		      end
		    default: NextState = S_0;                 
		    endcase
		    end
		end

	//--------------------------------------------------------------------------
endmodule
//------------------------------------------------------------------------------
