module Control(
  input   Clock,
  input   Reset,);
  //--|Parameters|--------------------------------------------------------------

  //--|Solution|----------------------------------------------------------------

endmodule
