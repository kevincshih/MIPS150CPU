module bios150v3(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c00043e;
30'h00000002: inst = 32'h37bd3000;
30'h00000003: inst = 32'h27bdffe0;
30'h00000004: inst = 32'h24020000;
30'h00000005: inst = 32'hafa40010;
30'h00000006: inst = 32'ha3a20014;
30'h00000007: inst = 32'hafa00018;
30'h00000008: inst = 32'h8fa20018;
30'h00000009: inst = 32'h00000000;
30'h0000000a: inst = 32'h2c420003;
30'h0000000b: inst = 32'h14400004;
30'h0000000c: inst = 32'h00000000;
30'h0000000d: inst = 32'h24020000;
30'h0000000e: inst = 32'h0800001a;
30'h0000000f: inst = 32'h00000000;
30'h00000010: inst = 32'h8fa20010;
30'h00000011: inst = 32'h00000000;
30'h00000012: inst = 32'h8fa30018;
30'h00000013: inst = 32'h00000000;
30'h00000014: inst = 32'h00431021;
30'h00000015: inst = 32'h80420000;
30'h00000016: inst = 32'h00000000;
30'h00000017: inst = 32'h24030000;
30'h00000018: inst = 32'h00431026;
30'h00000019: inst = 32'h0002102b;
30'h0000001a: inst = 32'h30420001;
30'h0000001b: inst = 32'h1040002b;
30'h0000001c: inst = 32'h00000000;
30'h0000001d: inst = 32'h8fa20010;
30'h0000001e: inst = 32'h00000000;
30'h0000001f: inst = 32'h8fa30018;
30'h00000020: inst = 32'h00000000;
30'h00000021: inst = 32'h00431021;
30'h00000022: inst = 32'h80420000;
30'h00000023: inst = 32'h00000000;
30'h00000024: inst = 32'h28420030;
30'h00000025: inst = 32'h1440001b;
30'h00000026: inst = 32'h00000000;
30'h00000027: inst = 32'h8fa20010;
30'h00000028: inst = 32'h00000000;
30'h00000029: inst = 32'h8fa30018;
30'h0000002a: inst = 32'h00000000;
30'h0000002b: inst = 32'h00431021;
30'h0000002c: inst = 32'h24030039;
30'h0000002d: inst = 32'h80420000;
30'h0000002e: inst = 32'h00000000;
30'h0000002f: inst = 32'h0062102a;
30'h00000030: inst = 32'h14400010;
30'h00000031: inst = 32'h00000000;
30'h00000032: inst = 32'h93a20014;
30'h00000033: inst = 32'h00000000;
30'h00000034: inst = 32'h8fa30018;
30'h00000035: inst = 32'h00000000;
30'h00000036: inst = 32'h8fa40010;
30'h00000037: inst = 32'h00000000;
30'h00000038: inst = 32'h00831821;
30'h00000039: inst = 32'h000220c0;
30'h0000003a: inst = 32'h00021040;
30'h0000003b: inst = 32'h90630000;
30'h0000003c: inst = 32'h00000000;
30'h0000003d: inst = 32'h00821021;
30'h0000003e: inst = 32'h00621021;
30'h0000003f: inst = 32'h2442ffd0;
30'h00000040: inst = 32'ha3a20014;
30'h00000041: inst = 32'h8fa20018;
30'h00000042: inst = 32'h00000000;
30'h00000043: inst = 32'h24420001;
30'h00000044: inst = 32'hafa20018;
30'h00000045: inst = 32'h08000008;
30'h00000046: inst = 32'h00000000;
30'h00000047: inst = 32'h93a20014;
30'h00000048: inst = 32'h00000000;
30'h00000049: inst = 32'h27bd0020;
30'h0000004a: inst = 32'h03e00008;
30'h0000004b: inst = 32'h00000000;
30'h0000004c: inst = 32'h27bdffe0;
30'h0000004d: inst = 32'h24020000;
30'h0000004e: inst = 32'hafa40010;
30'h0000004f: inst = 32'ha7a20014;
30'h00000050: inst = 32'hafa00018;
30'h00000051: inst = 32'h8fa20018;
30'h00000052: inst = 32'h00000000;
30'h00000053: inst = 32'h2c420005;
30'h00000054: inst = 32'h14400004;
30'h00000055: inst = 32'h00000000;
30'h00000056: inst = 32'h24020000;
30'h00000057: inst = 32'h08000063;
30'h00000058: inst = 32'h00000000;
30'h00000059: inst = 32'h8fa20010;
30'h0000005a: inst = 32'h00000000;
30'h0000005b: inst = 32'h8fa30018;
30'h0000005c: inst = 32'h00000000;
30'h0000005d: inst = 32'h00431021;
30'h0000005e: inst = 32'h80420000;
30'h0000005f: inst = 32'h00000000;
30'h00000060: inst = 32'h24030000;
30'h00000061: inst = 32'h00431026;
30'h00000062: inst = 32'h0002102b;
30'h00000063: inst = 32'h30420001;
30'h00000064: inst = 32'h1040002b;
30'h00000065: inst = 32'h00000000;
30'h00000066: inst = 32'h8fa20010;
30'h00000067: inst = 32'h00000000;
30'h00000068: inst = 32'h8fa30018;
30'h00000069: inst = 32'h00000000;
30'h0000006a: inst = 32'h00431021;
30'h0000006b: inst = 32'h80420000;
30'h0000006c: inst = 32'h00000000;
30'h0000006d: inst = 32'h28420030;
30'h0000006e: inst = 32'h1440001b;
30'h0000006f: inst = 32'h00000000;
30'h00000070: inst = 32'h8fa20010;
30'h00000071: inst = 32'h00000000;
30'h00000072: inst = 32'h8fa30018;
30'h00000073: inst = 32'h00000000;
30'h00000074: inst = 32'h00431021;
30'h00000075: inst = 32'h24030039;
30'h00000076: inst = 32'h80420000;
30'h00000077: inst = 32'h00000000;
30'h00000078: inst = 32'h0062102a;
30'h00000079: inst = 32'h14400010;
30'h0000007a: inst = 32'h00000000;
30'h0000007b: inst = 32'h97a20014;
30'h0000007c: inst = 32'h00000000;
30'h0000007d: inst = 32'h8fa30018;
30'h0000007e: inst = 32'h00000000;
30'h0000007f: inst = 32'h8fa40010;
30'h00000080: inst = 32'h00000000;
30'h00000081: inst = 32'h00831821;
30'h00000082: inst = 32'h000220c0;
30'h00000083: inst = 32'h00021040;
30'h00000084: inst = 32'h80630000;
30'h00000085: inst = 32'h00000000;
30'h00000086: inst = 32'h00821021;
30'h00000087: inst = 32'h00621021;
30'h00000088: inst = 32'h2442ffd0;
30'h00000089: inst = 32'ha7a20014;
30'h0000008a: inst = 32'h8fa20018;
30'h0000008b: inst = 32'h00000000;
30'h0000008c: inst = 32'h24420001;
30'h0000008d: inst = 32'hafa20018;
30'h0000008e: inst = 32'h08000051;
30'h0000008f: inst = 32'h00000000;
30'h00000090: inst = 32'h97a20014;
30'h00000091: inst = 32'h00000000;
30'h00000092: inst = 32'h27bd0020;
30'h00000093: inst = 32'h03e00008;
30'h00000094: inst = 32'h00000000;
30'h00000095: inst = 32'h27bdffe0;
30'h00000096: inst = 32'hafa40010;
30'h00000097: inst = 32'hafa00014;
30'h00000098: inst = 32'hafa00018;
30'h00000099: inst = 32'h8fa20018;
30'h0000009a: inst = 32'h00000000;
30'h0000009b: inst = 32'h2c420009;
30'h0000009c: inst = 32'h14400004;
30'h0000009d: inst = 32'h00000000;
30'h0000009e: inst = 32'h24020000;
30'h0000009f: inst = 32'h080000ab;
30'h000000a0: inst = 32'h00000000;
30'h000000a1: inst = 32'h8fa20010;
30'h000000a2: inst = 32'h00000000;
30'h000000a3: inst = 32'h8fa30018;
30'h000000a4: inst = 32'h00000000;
30'h000000a5: inst = 32'h00431021;
30'h000000a6: inst = 32'h80420000;
30'h000000a7: inst = 32'h00000000;
30'h000000a8: inst = 32'h24030000;
30'h000000a9: inst = 32'h00431026;
30'h000000aa: inst = 32'h0002102b;
30'h000000ab: inst = 32'h30420001;
30'h000000ac: inst = 32'h1040002b;
30'h000000ad: inst = 32'h00000000;
30'h000000ae: inst = 32'h8fa20010;
30'h000000af: inst = 32'h00000000;
30'h000000b0: inst = 32'h8fa30018;
30'h000000b1: inst = 32'h00000000;
30'h000000b2: inst = 32'h00431021;
30'h000000b3: inst = 32'h80420000;
30'h000000b4: inst = 32'h00000000;
30'h000000b5: inst = 32'h28420030;
30'h000000b6: inst = 32'h1440001b;
30'h000000b7: inst = 32'h00000000;
30'h000000b8: inst = 32'h8fa20010;
30'h000000b9: inst = 32'h00000000;
30'h000000ba: inst = 32'h8fa30018;
30'h000000bb: inst = 32'h00000000;
30'h000000bc: inst = 32'h00431021;
30'h000000bd: inst = 32'h24030039;
30'h000000be: inst = 32'h80420000;
30'h000000bf: inst = 32'h00000000;
30'h000000c0: inst = 32'h0062102a;
30'h000000c1: inst = 32'h14400010;
30'h000000c2: inst = 32'h00000000;
30'h000000c3: inst = 32'h8fa20014;
30'h000000c4: inst = 32'h00000000;
30'h000000c5: inst = 32'h8fa30018;
30'h000000c6: inst = 32'h00000000;
30'h000000c7: inst = 32'h8fa40010;
30'h000000c8: inst = 32'h00000000;
30'h000000c9: inst = 32'h00831821;
30'h000000ca: inst = 32'h000220c0;
30'h000000cb: inst = 32'h00021040;
30'h000000cc: inst = 32'h80630000;
30'h000000cd: inst = 32'h00000000;
30'h000000ce: inst = 32'h00821021;
30'h000000cf: inst = 32'h00621021;
30'h000000d0: inst = 32'h2442ffd0;
30'h000000d1: inst = 32'hafa20014;
30'h000000d2: inst = 32'h8fa20018;
30'h000000d3: inst = 32'h00000000;
30'h000000d4: inst = 32'h24420001;
30'h000000d5: inst = 32'hafa20018;
30'h000000d6: inst = 32'h08000099;
30'h000000d7: inst = 32'h00000000;
30'h000000d8: inst = 32'h8fa20014;
30'h000000d9: inst = 32'h00000000;
30'h000000da: inst = 32'h27bd0020;
30'h000000db: inst = 32'h03e00008;
30'h000000dc: inst = 32'h00000000;
30'h000000dd: inst = 32'h27bdffe0;
30'h000000de: inst = 32'h24020000;
30'h000000df: inst = 32'hafa40010;
30'h000000e0: inst = 32'ha3a20014;
30'h000000e1: inst = 32'ha3a20018;
30'h000000e2: inst = 32'h93a20018;
30'h000000e3: inst = 32'h00000000;
30'h000000e4: inst = 32'h2c420002;
30'h000000e5: inst = 32'h14400004;
30'h000000e6: inst = 32'h00000000;
30'h000000e7: inst = 32'h24020000;
30'h000000e8: inst = 32'h080000f4;
30'h000000e9: inst = 32'h00000000;
30'h000000ea: inst = 32'h8fa20010;
30'h000000eb: inst = 32'h00000000;
30'h000000ec: inst = 32'h93a30018;
30'h000000ed: inst = 32'h00000000;
30'h000000ee: inst = 32'h00431021;
30'h000000ef: inst = 32'h80420000;
30'h000000f0: inst = 32'h00000000;
30'h000000f1: inst = 32'h24030000;
30'h000000f2: inst = 32'h00431026;
30'h000000f3: inst = 32'h0002102b;
30'h000000f4: inst = 32'h30420001;
30'h000000f5: inst = 32'h1040006c;
30'h000000f6: inst = 32'h00000000;
30'h000000f7: inst = 32'h8fa20010;
30'h000000f8: inst = 32'h00000000;
30'h000000f9: inst = 32'h93a30018;
30'h000000fa: inst = 32'h00000000;
30'h000000fb: inst = 32'h00431021;
30'h000000fc: inst = 32'h80420000;
30'h000000fd: inst = 32'h00000000;
30'h000000fe: inst = 32'h28420030;
30'h000000ff: inst = 32'h14400019;
30'h00000100: inst = 32'h00000000;
30'h00000101: inst = 32'h8fa20010;
30'h00000102: inst = 32'h00000000;
30'h00000103: inst = 32'h93a30018;
30'h00000104: inst = 32'h00000000;
30'h00000105: inst = 32'h00431021;
30'h00000106: inst = 32'h24030039;
30'h00000107: inst = 32'h80420000;
30'h00000108: inst = 32'h00000000;
30'h00000109: inst = 32'h0062102a;
30'h0000010a: inst = 32'h1440000e;
30'h0000010b: inst = 32'h00000000;
30'h0000010c: inst = 32'h93a20018;
30'h0000010d: inst = 32'h00000000;
30'h0000010e: inst = 32'h8fa30010;
30'h0000010f: inst = 32'h00000000;
30'h00000110: inst = 32'h93a40014;
30'h00000111: inst = 32'h00000000;
30'h00000112: inst = 32'h00621021;
30'h00000113: inst = 32'h90420000;
30'h00000114: inst = 32'h00000000;
30'h00000115: inst = 32'h00041900;
30'h00000116: inst = 32'h00431021;
30'h00000117: inst = 32'h2442ffd0;
30'h00000118: inst = 32'ha3a20014;
30'h00000119: inst = 32'h8fa20010;
30'h0000011a: inst = 32'h00000000;
30'h0000011b: inst = 32'h93a30018;
30'h0000011c: inst = 32'h00000000;
30'h0000011d: inst = 32'h00431021;
30'h0000011e: inst = 32'h80420000;
30'h0000011f: inst = 32'h00000000;
30'h00000120: inst = 32'h28420061;
30'h00000121: inst = 32'h14400019;
30'h00000122: inst = 32'h00000000;
30'h00000123: inst = 32'h8fa20010;
30'h00000124: inst = 32'h00000000;
30'h00000125: inst = 32'h93a30018;
30'h00000126: inst = 32'h00000000;
30'h00000127: inst = 32'h00431021;
30'h00000128: inst = 32'h24030066;
30'h00000129: inst = 32'h80420000;
30'h0000012a: inst = 32'h00000000;
30'h0000012b: inst = 32'h0062102a;
30'h0000012c: inst = 32'h1440000e;
30'h0000012d: inst = 32'h00000000;
30'h0000012e: inst = 32'h93a20018;
30'h0000012f: inst = 32'h00000000;
30'h00000130: inst = 32'h8fa30010;
30'h00000131: inst = 32'h00000000;
30'h00000132: inst = 32'h93a40014;
30'h00000133: inst = 32'h00000000;
30'h00000134: inst = 32'h00621021;
30'h00000135: inst = 32'h90420000;
30'h00000136: inst = 32'h00000000;
30'h00000137: inst = 32'h00041900;
30'h00000138: inst = 32'h00431021;
30'h00000139: inst = 32'h2442ffa9;
30'h0000013a: inst = 32'ha3a20014;
30'h0000013b: inst = 32'h8fa20010;
30'h0000013c: inst = 32'h00000000;
30'h0000013d: inst = 32'h93a30018;
30'h0000013e: inst = 32'h00000000;
30'h0000013f: inst = 32'h00431021;
30'h00000140: inst = 32'h80420000;
30'h00000141: inst = 32'h00000000;
30'h00000142: inst = 32'h28420041;
30'h00000143: inst = 32'h14400019;
30'h00000144: inst = 32'h00000000;
30'h00000145: inst = 32'h8fa20010;
30'h00000146: inst = 32'h00000000;
30'h00000147: inst = 32'h93a30018;
30'h00000148: inst = 32'h00000000;
30'h00000149: inst = 32'h00431021;
30'h0000014a: inst = 32'h24030046;
30'h0000014b: inst = 32'h80420000;
30'h0000014c: inst = 32'h00000000;
30'h0000014d: inst = 32'h0062102a;
30'h0000014e: inst = 32'h1440000e;
30'h0000014f: inst = 32'h00000000;
30'h00000150: inst = 32'h93a20018;
30'h00000151: inst = 32'h00000000;
30'h00000152: inst = 32'h8fa30010;
30'h00000153: inst = 32'h00000000;
30'h00000154: inst = 32'h93a40014;
30'h00000155: inst = 32'h00000000;
30'h00000156: inst = 32'h00621021;
30'h00000157: inst = 32'h90420000;
30'h00000158: inst = 32'h00000000;
30'h00000159: inst = 32'h00041900;
30'h0000015a: inst = 32'h00431021;
30'h0000015b: inst = 32'h2442ffc9;
30'h0000015c: inst = 32'ha3a20014;
30'h0000015d: inst = 32'h93a20018;
30'h0000015e: inst = 32'h00000000;
30'h0000015f: inst = 32'h24420001;
30'h00000160: inst = 32'h080000e1;
30'h00000161: inst = 32'h00000000;
30'h00000162: inst = 32'h93a20014;
30'h00000163: inst = 32'h00000000;
30'h00000164: inst = 32'h27bd0020;
30'h00000165: inst = 32'h03e00008;
30'h00000166: inst = 32'h00000000;
30'h00000167: inst = 32'h27bdffe0;
30'h00000168: inst = 32'h24020000;
30'h00000169: inst = 32'hafa40010;
30'h0000016a: inst = 32'ha7a20014;
30'h0000016b: inst = 32'ha7a20018;
30'h0000016c: inst = 32'h97a20018;
30'h0000016d: inst = 32'h00000000;
30'h0000016e: inst = 32'h2c420004;
30'h0000016f: inst = 32'h14400004;
30'h00000170: inst = 32'h00000000;
30'h00000171: inst = 32'h24020000;
30'h00000172: inst = 32'h0800017e;
30'h00000173: inst = 32'h00000000;
30'h00000174: inst = 32'h8fa20010;
30'h00000175: inst = 32'h00000000;
30'h00000176: inst = 32'h97a30018;
30'h00000177: inst = 32'h00000000;
30'h00000178: inst = 32'h00431021;
30'h00000179: inst = 32'h80420000;
30'h0000017a: inst = 32'h00000000;
30'h0000017b: inst = 32'h24030000;
30'h0000017c: inst = 32'h00431026;
30'h0000017d: inst = 32'h0002102b;
30'h0000017e: inst = 32'h30420001;
30'h0000017f: inst = 32'h1040006c;
30'h00000180: inst = 32'h00000000;
30'h00000181: inst = 32'h8fa20010;
30'h00000182: inst = 32'h00000000;
30'h00000183: inst = 32'h97a30018;
30'h00000184: inst = 32'h00000000;
30'h00000185: inst = 32'h00431021;
30'h00000186: inst = 32'h80420000;
30'h00000187: inst = 32'h00000000;
30'h00000188: inst = 32'h28420030;
30'h00000189: inst = 32'h14400019;
30'h0000018a: inst = 32'h00000000;
30'h0000018b: inst = 32'h8fa20010;
30'h0000018c: inst = 32'h00000000;
30'h0000018d: inst = 32'h97a30018;
30'h0000018e: inst = 32'h00000000;
30'h0000018f: inst = 32'h00431021;
30'h00000190: inst = 32'h24030039;
30'h00000191: inst = 32'h80420000;
30'h00000192: inst = 32'h00000000;
30'h00000193: inst = 32'h0062102a;
30'h00000194: inst = 32'h1440000e;
30'h00000195: inst = 32'h00000000;
30'h00000196: inst = 32'h97a20018;
30'h00000197: inst = 32'h00000000;
30'h00000198: inst = 32'h8fa30010;
30'h00000199: inst = 32'h00000000;
30'h0000019a: inst = 32'h97a40014;
30'h0000019b: inst = 32'h00000000;
30'h0000019c: inst = 32'h00621021;
30'h0000019d: inst = 32'h80420000;
30'h0000019e: inst = 32'h00000000;
30'h0000019f: inst = 32'h00041900;
30'h000001a0: inst = 32'h00431021;
30'h000001a1: inst = 32'h2442ffd0;
30'h000001a2: inst = 32'ha7a20014;
30'h000001a3: inst = 32'h8fa20010;
30'h000001a4: inst = 32'h00000000;
30'h000001a5: inst = 32'h97a30018;
30'h000001a6: inst = 32'h00000000;
30'h000001a7: inst = 32'h00431021;
30'h000001a8: inst = 32'h80420000;
30'h000001a9: inst = 32'h00000000;
30'h000001aa: inst = 32'h28420061;
30'h000001ab: inst = 32'h14400019;
30'h000001ac: inst = 32'h00000000;
30'h000001ad: inst = 32'h8fa20010;
30'h000001ae: inst = 32'h00000000;
30'h000001af: inst = 32'h97a30018;
30'h000001b0: inst = 32'h00000000;
30'h000001b1: inst = 32'h00431021;
30'h000001b2: inst = 32'h24030066;
30'h000001b3: inst = 32'h80420000;
30'h000001b4: inst = 32'h00000000;
30'h000001b5: inst = 32'h0062102a;
30'h000001b6: inst = 32'h1440000e;
30'h000001b7: inst = 32'h00000000;
30'h000001b8: inst = 32'h97a20018;
30'h000001b9: inst = 32'h00000000;
30'h000001ba: inst = 32'h8fa30010;
30'h000001bb: inst = 32'h00000000;
30'h000001bc: inst = 32'h97a40014;
30'h000001bd: inst = 32'h00000000;
30'h000001be: inst = 32'h00621021;
30'h000001bf: inst = 32'h80420000;
30'h000001c0: inst = 32'h00000000;
30'h000001c1: inst = 32'h00041900;
30'h000001c2: inst = 32'h00431021;
30'h000001c3: inst = 32'h2442ffa9;
30'h000001c4: inst = 32'ha7a20014;
30'h000001c5: inst = 32'h8fa20010;
30'h000001c6: inst = 32'h00000000;
30'h000001c7: inst = 32'h97a30018;
30'h000001c8: inst = 32'h00000000;
30'h000001c9: inst = 32'h00431021;
30'h000001ca: inst = 32'h80420000;
30'h000001cb: inst = 32'h00000000;
30'h000001cc: inst = 32'h28420041;
30'h000001cd: inst = 32'h14400019;
30'h000001ce: inst = 32'h00000000;
30'h000001cf: inst = 32'h8fa20010;
30'h000001d0: inst = 32'h00000000;
30'h000001d1: inst = 32'h97a30018;
30'h000001d2: inst = 32'h00000000;
30'h000001d3: inst = 32'h00431021;
30'h000001d4: inst = 32'h24030046;
30'h000001d5: inst = 32'h80420000;
30'h000001d6: inst = 32'h00000000;
30'h000001d7: inst = 32'h0062102a;
30'h000001d8: inst = 32'h1440000e;
30'h000001d9: inst = 32'h00000000;
30'h000001da: inst = 32'h97a20018;
30'h000001db: inst = 32'h00000000;
30'h000001dc: inst = 32'h8fa30010;
30'h000001dd: inst = 32'h00000000;
30'h000001de: inst = 32'h97a40014;
30'h000001df: inst = 32'h00000000;
30'h000001e0: inst = 32'h00621021;
30'h000001e1: inst = 32'h80420000;
30'h000001e2: inst = 32'h00000000;
30'h000001e3: inst = 32'h00041900;
30'h000001e4: inst = 32'h00431021;
30'h000001e5: inst = 32'h2442ffc9;
30'h000001e6: inst = 32'ha7a20014;
30'h000001e7: inst = 32'h97a20018;
30'h000001e8: inst = 32'h00000000;
30'h000001e9: inst = 32'h24420001;
30'h000001ea: inst = 32'h0800016b;
30'h000001eb: inst = 32'h00000000;
30'h000001ec: inst = 32'h97a20014;
30'h000001ed: inst = 32'h00000000;
30'h000001ee: inst = 32'h27bd0020;
30'h000001ef: inst = 32'h03e00008;
30'h000001f0: inst = 32'h00000000;
30'h000001f1: inst = 32'h27bdffe0;
30'h000001f2: inst = 32'hafa40010;
30'h000001f3: inst = 32'hafa00014;
30'h000001f4: inst = 32'hafa00018;
30'h000001f5: inst = 32'h8fa20018;
30'h000001f6: inst = 32'h00000000;
30'h000001f7: inst = 32'h2c420008;
30'h000001f8: inst = 32'h14400004;
30'h000001f9: inst = 32'h00000000;
30'h000001fa: inst = 32'h24020000;
30'h000001fb: inst = 32'h08000207;
30'h000001fc: inst = 32'h00000000;
30'h000001fd: inst = 32'h8fa20010;
30'h000001fe: inst = 32'h00000000;
30'h000001ff: inst = 32'h8fa30018;
30'h00000200: inst = 32'h00000000;
30'h00000201: inst = 32'h00431021;
30'h00000202: inst = 32'h80420000;
30'h00000203: inst = 32'h00000000;
30'h00000204: inst = 32'h24030000;
30'h00000205: inst = 32'h00431026;
30'h00000206: inst = 32'h0002102b;
30'h00000207: inst = 32'h30420001;
30'h00000208: inst = 32'h1040006d;
30'h00000209: inst = 32'h00000000;
30'h0000020a: inst = 32'h8fa20010;
30'h0000020b: inst = 32'h00000000;
30'h0000020c: inst = 32'h8fa30018;
30'h0000020d: inst = 32'h00000000;
30'h0000020e: inst = 32'h00431021;
30'h0000020f: inst = 32'h80420000;
30'h00000210: inst = 32'h00000000;
30'h00000211: inst = 32'h28420030;
30'h00000212: inst = 32'h14400019;
30'h00000213: inst = 32'h00000000;
30'h00000214: inst = 32'h8fa20010;
30'h00000215: inst = 32'h00000000;
30'h00000216: inst = 32'h8fa30018;
30'h00000217: inst = 32'h00000000;
30'h00000218: inst = 32'h00431021;
30'h00000219: inst = 32'h24030039;
30'h0000021a: inst = 32'h80420000;
30'h0000021b: inst = 32'h00000000;
30'h0000021c: inst = 32'h0062102a;
30'h0000021d: inst = 32'h1440000e;
30'h0000021e: inst = 32'h00000000;
30'h0000021f: inst = 32'h8fa20018;
30'h00000220: inst = 32'h00000000;
30'h00000221: inst = 32'h8fa30010;
30'h00000222: inst = 32'h00000000;
30'h00000223: inst = 32'h8fa40014;
30'h00000224: inst = 32'h00000000;
30'h00000225: inst = 32'h00621021;
30'h00000226: inst = 32'h80420000;
30'h00000227: inst = 32'h00000000;
30'h00000228: inst = 32'h00041900;
30'h00000229: inst = 32'h00431021;
30'h0000022a: inst = 32'h2442ffd0;
30'h0000022b: inst = 32'hafa20014;
30'h0000022c: inst = 32'h8fa20010;
30'h0000022d: inst = 32'h00000000;
30'h0000022e: inst = 32'h8fa30018;
30'h0000022f: inst = 32'h00000000;
30'h00000230: inst = 32'h00431021;
30'h00000231: inst = 32'h80420000;
30'h00000232: inst = 32'h00000000;
30'h00000233: inst = 32'h28420061;
30'h00000234: inst = 32'h14400019;
30'h00000235: inst = 32'h00000000;
30'h00000236: inst = 32'h8fa20010;
30'h00000237: inst = 32'h00000000;
30'h00000238: inst = 32'h8fa30018;
30'h00000239: inst = 32'h00000000;
30'h0000023a: inst = 32'h00431021;
30'h0000023b: inst = 32'h24030066;
30'h0000023c: inst = 32'h80420000;
30'h0000023d: inst = 32'h00000000;
30'h0000023e: inst = 32'h0062102a;
30'h0000023f: inst = 32'h1440000e;
30'h00000240: inst = 32'h00000000;
30'h00000241: inst = 32'h8fa20018;
30'h00000242: inst = 32'h00000000;
30'h00000243: inst = 32'h8fa30010;
30'h00000244: inst = 32'h00000000;
30'h00000245: inst = 32'h8fa40014;
30'h00000246: inst = 32'h00000000;
30'h00000247: inst = 32'h00621021;
30'h00000248: inst = 32'h80420000;
30'h00000249: inst = 32'h00000000;
30'h0000024a: inst = 32'h00041900;
30'h0000024b: inst = 32'h00431021;
30'h0000024c: inst = 32'h2442ffa9;
30'h0000024d: inst = 32'hafa20014;
30'h0000024e: inst = 32'h8fa20010;
30'h0000024f: inst = 32'h00000000;
30'h00000250: inst = 32'h8fa30018;
30'h00000251: inst = 32'h00000000;
30'h00000252: inst = 32'h00431021;
30'h00000253: inst = 32'h80420000;
30'h00000254: inst = 32'h00000000;
30'h00000255: inst = 32'h28420041;
30'h00000256: inst = 32'h14400019;
30'h00000257: inst = 32'h00000000;
30'h00000258: inst = 32'h8fa20010;
30'h00000259: inst = 32'h00000000;
30'h0000025a: inst = 32'h8fa30018;
30'h0000025b: inst = 32'h00000000;
30'h0000025c: inst = 32'h00431021;
30'h0000025d: inst = 32'h24030046;
30'h0000025e: inst = 32'h80420000;
30'h0000025f: inst = 32'h00000000;
30'h00000260: inst = 32'h0062102a;
30'h00000261: inst = 32'h1440000e;
30'h00000262: inst = 32'h00000000;
30'h00000263: inst = 32'h8fa20018;
30'h00000264: inst = 32'h00000000;
30'h00000265: inst = 32'h8fa30010;
30'h00000266: inst = 32'h00000000;
30'h00000267: inst = 32'h8fa40014;
30'h00000268: inst = 32'h00000000;
30'h00000269: inst = 32'h00621021;
30'h0000026a: inst = 32'h80420000;
30'h0000026b: inst = 32'h00000000;
30'h0000026c: inst = 32'h00041900;
30'h0000026d: inst = 32'h00431021;
30'h0000026e: inst = 32'h2442ffc9;
30'h0000026f: inst = 32'hafa20014;
30'h00000270: inst = 32'h8fa20018;
30'h00000271: inst = 32'h00000000;
30'h00000272: inst = 32'h24420001;
30'h00000273: inst = 32'hafa20018;
30'h00000274: inst = 32'h080001f5;
30'h00000275: inst = 32'h00000000;
30'h00000276: inst = 32'h8fa20014;
30'h00000277: inst = 32'h00000000;
30'h00000278: inst = 32'h27bd0020;
30'h00000279: inst = 32'h03e00008;
30'h0000027a: inst = 32'h00000000;
30'h0000027b: inst = 32'h27bdffd8;
30'h0000027c: inst = 32'ha3a40010;
30'h0000027d: inst = 32'hafa50014;
30'h0000027e: inst = 32'hafa60018;
30'h0000027f: inst = 32'h24020002;
30'h00000280: inst = 32'hafa0001c;
30'h00000281: inst = 32'hafa20020;
30'h00000282: inst = 32'h8fa2001c;
30'h00000283: inst = 32'h00000000;
30'h00000284: inst = 32'h8fa30020;
30'h00000285: inst = 32'h00000000;
30'h00000286: inst = 32'h0043102b;
30'h00000287: inst = 32'h14400004;
30'h00000288: inst = 32'h00000000;
30'h00000289: inst = 32'h24020000;
30'h0000028a: inst = 32'h08000292;
30'h0000028b: inst = 32'h00000000;
30'h0000028c: inst = 32'h8fa2001c;
30'h0000028d: inst = 32'h00000000;
30'h0000028e: inst = 32'h24420001;
30'h0000028f: inst = 32'h8fa30018;
30'h00000290: inst = 32'h00000000;
30'h00000291: inst = 32'h0043102b;
30'h00000292: inst = 32'h30420001;
30'h00000293: inst = 32'h1040003a;
30'h00000294: inst = 32'h00000000;
30'h00000295: inst = 32'h8fa20020;
30'h00000296: inst = 32'h00000000;
30'h00000297: inst = 32'h2442ffff;
30'h00000298: inst = 32'h8fa3001c;
30'h00000299: inst = 32'h00000000;
30'h0000029a: inst = 32'h00431023;
30'h0000029b: inst = 32'h93a30010;
30'h0000029c: inst = 32'h00000000;
30'h0000029d: inst = 32'h00021080;
30'h0000029e: inst = 32'h00431006;
30'h0000029f: inst = 32'h3042000f;
30'h000002a0: inst = 32'ha3a20024;
30'h000002a1: inst = 32'h83a20024;
30'h000002a2: inst = 32'h00000000;
30'h000002a3: inst = 32'h04400010;
30'h000002a4: inst = 32'h00000000;
30'h000002a5: inst = 32'h24020009;
30'h000002a6: inst = 32'h83a30024;
30'h000002a7: inst = 32'h00000000;
30'h000002a8: inst = 32'h0043102a;
30'h000002a9: inst = 32'h1440000a;
30'h000002aa: inst = 32'h00000000;
30'h000002ab: inst = 32'h93a20024;
30'h000002ac: inst = 32'h00000000;
30'h000002ad: inst = 32'h8fa3001c;
30'h000002ae: inst = 32'h00000000;
30'h000002af: inst = 32'h8fa40014;
30'h000002b0: inst = 32'h00000000;
30'h000002b1: inst = 32'h24420030;
30'h000002b2: inst = 32'h00831821;
30'h000002b3: inst = 32'ha0620000;
30'h000002b4: inst = 32'h83a20024;
30'h000002b5: inst = 32'h00000000;
30'h000002b6: inst = 32'h2842000a;
30'h000002b7: inst = 32'h14400010;
30'h000002b8: inst = 32'h00000000;
30'h000002b9: inst = 32'h2402000f;
30'h000002ba: inst = 32'h83a30024;
30'h000002bb: inst = 32'h00000000;
30'h000002bc: inst = 32'h0043102a;
30'h000002bd: inst = 32'h1440000a;
30'h000002be: inst = 32'h00000000;
30'h000002bf: inst = 32'h93a20024;
30'h000002c0: inst = 32'h00000000;
30'h000002c1: inst = 32'h8fa3001c;
30'h000002c2: inst = 32'h00000000;
30'h000002c3: inst = 32'h8fa40014;
30'h000002c4: inst = 32'h00000000;
30'h000002c5: inst = 32'h24420057;
30'h000002c6: inst = 32'h00831821;
30'h000002c7: inst = 32'ha0620000;
30'h000002c8: inst = 32'h8fa2001c;
30'h000002c9: inst = 32'h00000000;
30'h000002ca: inst = 32'h24420001;
30'h000002cb: inst = 32'hafa2001c;
30'h000002cc: inst = 32'h08000282;
30'h000002cd: inst = 32'h00000000;
30'h000002ce: inst = 32'h8fa2001c;
30'h000002cf: inst = 32'h00000000;
30'h000002d0: inst = 32'h8fa30014;
30'h000002d1: inst = 32'h00000000;
30'h000002d2: inst = 32'h24040000;
30'h000002d3: inst = 32'h00621021;
30'h000002d4: inst = 32'ha0440000;
30'h000002d5: inst = 32'h8fa20014;
30'h000002d6: inst = 32'h00000000;
30'h000002d7: inst = 32'h27bd0028;
30'h000002d8: inst = 32'h03e00008;
30'h000002d9: inst = 32'h00000000;
30'h000002da: inst = 32'h27bdffd8;
30'h000002db: inst = 32'ha7a40010;
30'h000002dc: inst = 32'hafa50014;
30'h000002dd: inst = 32'hafa60018;
30'h000002de: inst = 32'h24020004;
30'h000002df: inst = 32'hafa0001c;
30'h000002e0: inst = 32'hafa20020;
30'h000002e1: inst = 32'h8fa2001c;
30'h000002e2: inst = 32'h00000000;
30'h000002e3: inst = 32'h8fa30020;
30'h000002e4: inst = 32'h00000000;
30'h000002e5: inst = 32'h0043102b;
30'h000002e6: inst = 32'h14400004;
30'h000002e7: inst = 32'h00000000;
30'h000002e8: inst = 32'h24020000;
30'h000002e9: inst = 32'h080002f1;
30'h000002ea: inst = 32'h00000000;
30'h000002eb: inst = 32'h8fa2001c;
30'h000002ec: inst = 32'h00000000;
30'h000002ed: inst = 32'h24420001;
30'h000002ee: inst = 32'h8fa30018;
30'h000002ef: inst = 32'h00000000;
30'h000002f0: inst = 32'h0043102b;
30'h000002f1: inst = 32'h30420001;
30'h000002f2: inst = 32'h1040003a;
30'h000002f3: inst = 32'h00000000;
30'h000002f4: inst = 32'h8fa20020;
30'h000002f5: inst = 32'h00000000;
30'h000002f6: inst = 32'h2442ffff;
30'h000002f7: inst = 32'h8fa3001c;
30'h000002f8: inst = 32'h00000000;
30'h000002f9: inst = 32'h00431023;
30'h000002fa: inst = 32'h97a30010;
30'h000002fb: inst = 32'h00000000;
30'h000002fc: inst = 32'h00021080;
30'h000002fd: inst = 32'h00431006;
30'h000002fe: inst = 32'h3042000f;
30'h000002ff: inst = 32'ha3a20024;
30'h00000300: inst = 32'h83a20024;
30'h00000301: inst = 32'h00000000;
30'h00000302: inst = 32'h04400010;
30'h00000303: inst = 32'h00000000;
30'h00000304: inst = 32'h24020009;
30'h00000305: inst = 32'h83a30024;
30'h00000306: inst = 32'h00000000;
30'h00000307: inst = 32'h0043102a;
30'h00000308: inst = 32'h1440000a;
30'h00000309: inst = 32'h00000000;
30'h0000030a: inst = 32'h93a20024;
30'h0000030b: inst = 32'h00000000;
30'h0000030c: inst = 32'h8fa3001c;
30'h0000030d: inst = 32'h00000000;
30'h0000030e: inst = 32'h8fa40014;
30'h0000030f: inst = 32'h00000000;
30'h00000310: inst = 32'h24420030;
30'h00000311: inst = 32'h00831821;
30'h00000312: inst = 32'ha0620000;
30'h00000313: inst = 32'h83a20024;
30'h00000314: inst = 32'h00000000;
30'h00000315: inst = 32'h2842000a;
30'h00000316: inst = 32'h14400010;
30'h00000317: inst = 32'h00000000;
30'h00000318: inst = 32'h2402000f;
30'h00000319: inst = 32'h83a30024;
30'h0000031a: inst = 32'h00000000;
30'h0000031b: inst = 32'h0043102a;
30'h0000031c: inst = 32'h1440000a;
30'h0000031d: inst = 32'h00000000;
30'h0000031e: inst = 32'h93a20024;
30'h0000031f: inst = 32'h00000000;
30'h00000320: inst = 32'h8fa3001c;
30'h00000321: inst = 32'h00000000;
30'h00000322: inst = 32'h8fa40014;
30'h00000323: inst = 32'h00000000;
30'h00000324: inst = 32'h24420057;
30'h00000325: inst = 32'h00831821;
30'h00000326: inst = 32'ha0620000;
30'h00000327: inst = 32'h8fa2001c;
30'h00000328: inst = 32'h00000000;
30'h00000329: inst = 32'h24420001;
30'h0000032a: inst = 32'hafa2001c;
30'h0000032b: inst = 32'h080002e1;
30'h0000032c: inst = 32'h00000000;
30'h0000032d: inst = 32'h8fa2001c;
30'h0000032e: inst = 32'h00000000;
30'h0000032f: inst = 32'h8fa30014;
30'h00000330: inst = 32'h00000000;
30'h00000331: inst = 32'h24040000;
30'h00000332: inst = 32'h00621021;
30'h00000333: inst = 32'ha0440000;
30'h00000334: inst = 32'h8fa20014;
30'h00000335: inst = 32'h00000000;
30'h00000336: inst = 32'h27bd0028;
30'h00000337: inst = 32'h03e00008;
30'h00000338: inst = 32'h00000000;
30'h00000339: inst = 32'h27bdffd8;
30'h0000033a: inst = 32'hafa40010;
30'h0000033b: inst = 32'hafa50014;
30'h0000033c: inst = 32'hafa60018;
30'h0000033d: inst = 32'h24020008;
30'h0000033e: inst = 32'hafa0001c;
30'h0000033f: inst = 32'hafa20020;
30'h00000340: inst = 32'h8fa2001c;
30'h00000341: inst = 32'h00000000;
30'h00000342: inst = 32'h8fa30020;
30'h00000343: inst = 32'h00000000;
30'h00000344: inst = 32'h0043102b;
30'h00000345: inst = 32'h14400004;
30'h00000346: inst = 32'h00000000;
30'h00000347: inst = 32'h24020000;
30'h00000348: inst = 32'h08000350;
30'h00000349: inst = 32'h00000000;
30'h0000034a: inst = 32'h8fa2001c;
30'h0000034b: inst = 32'h00000000;
30'h0000034c: inst = 32'h24420001;
30'h0000034d: inst = 32'h8fa30018;
30'h0000034e: inst = 32'h00000000;
30'h0000034f: inst = 32'h0043102b;
30'h00000350: inst = 32'h30420001;
30'h00000351: inst = 32'h1040003a;
30'h00000352: inst = 32'h00000000;
30'h00000353: inst = 32'h8fa20020;
30'h00000354: inst = 32'h00000000;
30'h00000355: inst = 32'h2442ffff;
30'h00000356: inst = 32'h8fa3001c;
30'h00000357: inst = 32'h00000000;
30'h00000358: inst = 32'h00431023;
30'h00000359: inst = 32'h8fa30010;
30'h0000035a: inst = 32'h00000000;
30'h0000035b: inst = 32'h00021080;
30'h0000035c: inst = 32'h00431006;
30'h0000035d: inst = 32'h3042000f;
30'h0000035e: inst = 32'ha3a20024;
30'h0000035f: inst = 32'h83a20024;
30'h00000360: inst = 32'h00000000;
30'h00000361: inst = 32'h04400010;
30'h00000362: inst = 32'h00000000;
30'h00000363: inst = 32'h24020009;
30'h00000364: inst = 32'h83a30024;
30'h00000365: inst = 32'h00000000;
30'h00000366: inst = 32'h0043102a;
30'h00000367: inst = 32'h1440000a;
30'h00000368: inst = 32'h00000000;
30'h00000369: inst = 32'h93a20024;
30'h0000036a: inst = 32'h00000000;
30'h0000036b: inst = 32'h8fa3001c;
30'h0000036c: inst = 32'h00000000;
30'h0000036d: inst = 32'h8fa40014;
30'h0000036e: inst = 32'h00000000;
30'h0000036f: inst = 32'h24420030;
30'h00000370: inst = 32'h00831821;
30'h00000371: inst = 32'ha0620000;
30'h00000372: inst = 32'h83a20024;
30'h00000373: inst = 32'h00000000;
30'h00000374: inst = 32'h2842000a;
30'h00000375: inst = 32'h14400010;
30'h00000376: inst = 32'h00000000;
30'h00000377: inst = 32'h2402000f;
30'h00000378: inst = 32'h83a30024;
30'h00000379: inst = 32'h00000000;
30'h0000037a: inst = 32'h0043102a;
30'h0000037b: inst = 32'h1440000a;
30'h0000037c: inst = 32'h00000000;
30'h0000037d: inst = 32'h93a20024;
30'h0000037e: inst = 32'h00000000;
30'h0000037f: inst = 32'h8fa3001c;
30'h00000380: inst = 32'h00000000;
30'h00000381: inst = 32'h8fa40014;
30'h00000382: inst = 32'h00000000;
30'h00000383: inst = 32'h24420057;
30'h00000384: inst = 32'h00831821;
30'h00000385: inst = 32'ha0620000;
30'h00000386: inst = 32'h8fa2001c;
30'h00000387: inst = 32'h00000000;
30'h00000388: inst = 32'h24420001;
30'h00000389: inst = 32'hafa2001c;
30'h0000038a: inst = 32'h08000340;
30'h0000038b: inst = 32'h00000000;
30'h0000038c: inst = 32'h8fa2001c;
30'h0000038d: inst = 32'h00000000;
30'h0000038e: inst = 32'h8fa30014;
30'h0000038f: inst = 32'h00000000;
30'h00000390: inst = 32'h24040000;
30'h00000391: inst = 32'h00621021;
30'h00000392: inst = 32'ha0440000;
30'h00000393: inst = 32'h8fa20014;
30'h00000394: inst = 32'h00000000;
30'h00000395: inst = 32'h27bd0028;
30'h00000396: inst = 32'h03e00008;
30'h00000397: inst = 32'h00000000;
30'h00000398: inst = 32'h27bdffc8;
30'h00000399: inst = 32'hafbf0034;
30'h0000039a: inst = 32'hafa40020;
30'h0000039b: inst = 32'hafa50024;
30'h0000039c: inst = 32'hafa00028;
30'h0000039d: inst = 32'h8fa20028;
30'h0000039e: inst = 32'h00000000;
30'h0000039f: inst = 32'h8fa30024;
30'h000003a0: inst = 32'h00000000;
30'h000003a1: inst = 32'h0043102b;
30'h000003a2: inst = 32'h1040000f;
30'h000003a3: inst = 32'h00000000;
30'h000003a4: inst = 32'h0c000635;
30'h000003a5: inst = 32'h00000000;
30'h000003a6: inst = 32'h8fa30028;
30'h000003a7: inst = 32'h00000000;
30'h000003a8: inst = 32'h8fa40020;
30'h000003a9: inst = 32'h00000000;
30'h000003aa: inst = 32'h00831821;
30'h000003ab: inst = 32'ha0620000;
30'h000003ac: inst = 32'h8fa20028;
30'h000003ad: inst = 32'h00000000;
30'h000003ae: inst = 32'h24420001;
30'h000003af: inst = 32'hafa20028;
30'h000003b0: inst = 32'h0800039d;
30'h000003b1: inst = 32'h00000000;
30'h000003b2: inst = 32'h8fa20024;
30'h000003b3: inst = 32'h00000000;
30'h000003b4: inst = 32'h8fa30020;
30'h000003b5: inst = 32'h00000000;
30'h000003b6: inst = 32'h24040000;
30'h000003b7: inst = 32'h00621021;
30'h000003b8: inst = 32'ha0440000;
30'h000003b9: inst = 32'h8fa20020;
30'h000003ba: inst = 32'h00000000;
30'h000003bb: inst = 32'h8fbf0034;
30'h000003bc: inst = 32'h00000000;
30'h000003bd: inst = 32'h27bd0038;
30'h000003be: inst = 32'h03e00008;
30'h000003bf: inst = 32'h00000000;
30'h000003c0: inst = 32'h27bdffb8;
30'h000003c1: inst = 32'hafbf0044;
30'h000003c2: inst = 32'hafa40024;
30'h000003c3: inst = 32'hafa50028;
30'h000003c4: inst = 32'hafa6002c;
30'h000003c5: inst = 32'hafa00030;
30'h000003c6: inst = 32'h8fa20030;
30'h000003c7: inst = 32'h00000000;
30'h000003c8: inst = 32'h8fa30028;
30'h000003c9: inst = 32'h00000000;
30'h000003ca: inst = 32'h0043102b;
30'h000003cb: inst = 32'h10400036;
30'h000003cc: inst = 32'h00000000;
30'h000003cd: inst = 32'h0c000635;
30'h000003ce: inst = 32'h00000000;
30'h000003cf: inst = 32'ha3a20034;
30'h000003d0: inst = 32'hafa00038;
30'h000003d1: inst = 32'h8fa2002c;
30'h000003d2: inst = 32'h00000000;
30'h000003d3: inst = 32'h8fa30038;
30'h000003d4: inst = 32'h00000000;
30'h000003d5: inst = 32'h00431021;
30'h000003d6: inst = 32'h80420000;
30'h000003d7: inst = 32'h00000000;
30'h000003d8: inst = 32'h1040001b;
30'h000003d9: inst = 32'h00000000;
30'h000003da: inst = 32'h8fa2002c;
30'h000003db: inst = 32'h00000000;
30'h000003dc: inst = 32'h8fa30038;
30'h000003dd: inst = 32'h00000000;
30'h000003de: inst = 32'h00431021;
30'h000003df: inst = 32'h83a30034;
30'h000003e0: inst = 32'h00000000;
30'h000003e1: inst = 32'h80420000;
30'h000003e2: inst = 32'h00000000;
30'h000003e3: inst = 32'h1462000a;
30'h000003e4: inst = 32'h00000000;
30'h000003e5: inst = 32'h8fa20030;
30'h000003e6: inst = 32'h00000000;
30'h000003e7: inst = 32'h8fa30024;
30'h000003e8: inst = 32'h00000000;
30'h000003e9: inst = 32'h24040000;
30'h000003ea: inst = 32'h00621021;
30'h000003eb: inst = 32'ha0440000;
30'h000003ec: inst = 32'h08000409;
30'h000003ed: inst = 32'h00000000;
30'h000003ee: inst = 32'h8fa20038;
30'h000003ef: inst = 32'h00000000;
30'h000003f0: inst = 32'h24420001;
30'h000003f1: inst = 32'hafa20038;
30'h000003f2: inst = 32'h080003d1;
30'h000003f3: inst = 32'h00000000;
30'h000003f4: inst = 32'h93a20034;
30'h000003f5: inst = 32'h00000000;
30'h000003f6: inst = 32'h8fa30030;
30'h000003f7: inst = 32'h00000000;
30'h000003f8: inst = 32'h8fa40024;
30'h000003f9: inst = 32'h00000000;
30'h000003fa: inst = 32'h00831821;
30'h000003fb: inst = 32'ha0620000;
30'h000003fc: inst = 32'h8fa20030;
30'h000003fd: inst = 32'h00000000;
30'h000003fe: inst = 32'h24420001;
30'h000003ff: inst = 32'hafa20030;
30'h00000400: inst = 32'h080003c6;
30'h00000401: inst = 32'h00000000;
30'h00000402: inst = 32'h8fa20028;
30'h00000403: inst = 32'h00000000;
30'h00000404: inst = 32'h8fa30024;
30'h00000405: inst = 32'h00000000;
30'h00000406: inst = 32'h24040000;
30'h00000407: inst = 32'h00431021;
30'h00000408: inst = 32'ha044ffff;
30'h00000409: inst = 32'h8fa20024;
30'h0000040a: inst = 32'h00000000;
30'h0000040b: inst = 32'hafa20020;
30'h0000040c: inst = 32'h8fa20020;
30'h0000040d: inst = 32'h00000000;
30'h0000040e: inst = 32'h8fbf0044;
30'h0000040f: inst = 32'h00000000;
30'h00000410: inst = 32'h27bd0048;
30'h00000411: inst = 32'h03e00008;
30'h00000412: inst = 32'h00000000;
30'h00000413: inst = 32'h27bdffb8;
30'h00000414: inst = 32'hafbf0044;
30'h00000415: inst = 32'hafa40020;
30'h00000416: inst = 32'hafa50024;
30'h00000417: inst = 32'hafa00028;
30'h00000418: inst = 32'h8fa20028;
30'h00000419: inst = 32'h00000000;
30'h0000041a: inst = 32'h00021080;
30'h0000041b: inst = 32'h8fa30024;
30'h0000041c: inst = 32'h00000000;
30'h0000041d: inst = 32'h0043102b;
30'h0000041e: inst = 32'h1040001a;
30'h0000041f: inst = 32'h00000000;
30'h00000420: inst = 32'h27a4002c;
30'h00000421: inst = 32'h24050008;
30'h00000422: inst = 32'h0c000398;
30'h00000423: inst = 32'h00000000;
30'h00000424: inst = 32'hafa20038;
30'h00000425: inst = 32'h8fa20028;
30'h00000426: inst = 32'h00000000;
30'h00000427: inst = 32'h8fa30020;
30'h00000428: inst = 32'h00000000;
30'h00000429: inst = 32'h00021080;
30'h0000042a: inst = 32'h00621021;
30'h0000042b: inst = 32'hafa2003c;
30'h0000042c: inst = 32'h8fa40038;
30'h0000042d: inst = 32'h00000000;
30'h0000042e: inst = 32'h0c0001f1;
30'h0000042f: inst = 32'h00000000;
30'h00000430: inst = 32'h8fa3003c;
30'h00000431: inst = 32'h00000000;
30'h00000432: inst = 32'hac620000;
30'h00000433: inst = 32'h8fa20028;
30'h00000434: inst = 32'h00000000;
30'h00000435: inst = 32'h24420001;
30'h00000436: inst = 32'hafa20028;
30'h00000437: inst = 32'h08000418;
30'h00000438: inst = 32'h00000000;
30'h00000439: inst = 32'h8fbf0044;
30'h0000043a: inst = 32'h00000000;
30'h0000043b: inst = 32'h27bd0048;
30'h0000043c: inst = 32'h03e00008;
30'h0000043d: inst = 32'h00000000;
30'h0000043e: inst = 32'h27bdfef0;
30'h0000043f: inst = 32'hafbf0108;
30'h00000440: inst = 32'hafb000f8;
30'h00000441: inst = 32'hafb100fc;
30'h00000442: inst = 32'hafb20100;
30'h00000443: inst = 32'hafa00020;
30'h00000444: inst = 32'h3c021000;
30'h00000445: inst = 32'h24441964;
30'h00000446: inst = 32'h0c000614;
30'h00000447: inst = 32'h00000000;
30'h00000448: inst = 32'h3c021000;
30'h00000449: inst = 32'h24441970;
30'h0000044a: inst = 32'h0c000614;
30'h0000044b: inst = 32'h00000000;
30'h0000044c: inst = 32'h3c021000;
30'h0000044d: inst = 32'h27a40024;
30'h0000044e: inst = 32'h24050080;
30'h0000044f: inst = 32'h24461974;
30'h00000450: inst = 32'h0c0003c0;
30'h00000451: inst = 32'h00000000;
30'h00000452: inst = 32'hafa200a4;
30'h00000453: inst = 32'h3c031000;
30'h00000454: inst = 32'h24651978;
30'h00000455: inst = 32'h00022021;
30'h00000456: inst = 32'h0c0005c1;
30'h00000457: inst = 32'h00000000;
30'h00000458: inst = 32'h1440001e;
30'h00000459: inst = 32'h00000000;
30'h0000045a: inst = 32'h3c021000;
30'h0000045b: inst = 32'h27b00024;
30'h0000045c: inst = 32'h24110080;
30'h0000045d: inst = 32'h24521974;
30'h0000045e: inst = 32'h00102021;
30'h0000045f: inst = 32'h00112821;
30'h00000460: inst = 32'h00123021;
30'h00000461: inst = 32'h0c0003c0;
30'h00000462: inst = 32'h00000000;
30'h00000463: inst = 32'h00022021;
30'h00000464: inst = 32'h0c0001f1;
30'h00000465: inst = 32'h00000000;
30'h00000466: inst = 32'hafa200a8;
30'h00000467: inst = 32'h00102021;
30'h00000468: inst = 32'h00112821;
30'h00000469: inst = 32'h00123021;
30'h0000046a: inst = 32'h0c0003c0;
30'h0000046b: inst = 32'h00000000;
30'h0000046c: inst = 32'h00022021;
30'h0000046d: inst = 32'h0c000095;
30'h0000046e: inst = 32'h00000000;
30'h0000046f: inst = 32'hafa200ac;
30'h00000470: inst = 32'h8fa400a8;
30'h00000471: inst = 32'h00000000;
30'h00000472: inst = 32'h00022821;
30'h00000473: inst = 32'h0c000413;
30'h00000474: inst = 32'h00000000;
30'h00000475: inst = 32'h08000448;
30'h00000476: inst = 32'h00000000;
30'h00000477: inst = 32'h8fa400a4;
30'h00000478: inst = 32'h00000000;
30'h00000479: inst = 32'h3c021000;
30'h0000047a: inst = 32'h24451980;
30'h0000047b: inst = 32'h0c0005c1;
30'h0000047c: inst = 32'h00000000;
30'h0000047d: inst = 32'h14400010;
30'h0000047e: inst = 32'h00000000;
30'h0000047f: inst = 32'h3c021000;
30'h00000480: inst = 32'h27a40024;
30'h00000481: inst = 32'h24050080;
30'h00000482: inst = 32'h24461974;
30'h00000483: inst = 32'h0c0003c0;
30'h00000484: inst = 32'h00000000;
30'h00000485: inst = 32'h00022021;
30'h00000486: inst = 32'h0c0001f1;
30'h00000487: inst = 32'h00000000;
30'h00000488: inst = 32'hafa200b0;
30'h00000489: inst = 32'hafa200b4;
30'h0000048a: inst = 32'h0040f809;
30'h0000048b: inst = 32'h00000000;
30'h0000048c: inst = 32'h08000448;
30'h0000048d: inst = 32'h00000000;
30'h0000048e: inst = 32'h8fa400a4;
30'h0000048f: inst = 32'h00000000;
30'h00000490: inst = 32'h3c021000;
30'h00000491: inst = 32'h24451984;
30'h00000492: inst = 32'h0c0005c1;
30'h00000493: inst = 32'h00000000;
30'h00000494: inst = 32'h1440002a;
30'h00000495: inst = 32'h00000000;
30'h00000496: inst = 32'h3c021000;
30'h00000497: inst = 32'h24461974;
30'h00000498: inst = 32'h27b00024;
30'h00000499: inst = 32'h24110080;
30'h0000049a: inst = 32'h00102021;
30'h0000049b: inst = 32'h00112821;
30'h0000049c: inst = 32'h0c0003c0;
30'h0000049d: inst = 32'h00000000;
30'h0000049e: inst = 32'h00022021;
30'h0000049f: inst = 32'h0c0001f1;
30'h000004a0: inst = 32'h00000000;
30'h000004a1: inst = 32'hafa200b8;
30'h000004a2: inst = 32'hafa200bc;
30'h000004a3: inst = 32'h8fa400b8;
30'h000004a4: inst = 32'h00000000;
30'h000004a5: inst = 32'h00102821;
30'h000004a6: inst = 32'h00113021;
30'h000004a7: inst = 32'h0c000339;
30'h000004a8: inst = 32'h00000000;
30'h000004a9: inst = 32'h00022021;
30'h000004aa: inst = 32'h0c000614;
30'h000004ab: inst = 32'h00000000;
30'h000004ac: inst = 32'h3c021000;
30'h000004ad: inst = 32'h24441988;
30'h000004ae: inst = 32'h0c000614;
30'h000004af: inst = 32'h00000000;
30'h000004b0: inst = 32'h8fa200bc;
30'h000004b1: inst = 32'h00000000;
30'h000004b2: inst = 32'h8c440000;
30'h000004b3: inst = 32'h00000000;
30'h000004b4: inst = 32'h00102821;
30'h000004b5: inst = 32'h00113021;
30'h000004b6: inst = 32'h0c000339;
30'h000004b7: inst = 32'h00000000;
30'h000004b8: inst = 32'h00022021;
30'h000004b9: inst = 32'h0c000614;
30'h000004ba: inst = 32'h00000000;
30'h000004bb: inst = 32'h3c021000;
30'h000004bc: inst = 32'h2444198c;
30'h000004bd: inst = 32'h08000446;
30'h000004be: inst = 32'h00000000;
30'h000004bf: inst = 32'h8fa400a4;
30'h000004c0: inst = 32'h00000000;
30'h000004c1: inst = 32'h3c021000;
30'h000004c2: inst = 32'h24451990;
30'h000004c3: inst = 32'h0c0005c1;
30'h000004c4: inst = 32'h00000000;
30'h000004c5: inst = 32'h14400025;
30'h000004c6: inst = 32'h00000000;
30'h000004c7: inst = 32'h3c021000;
30'h000004c8: inst = 32'h24461974;
30'h000004c9: inst = 32'h27b00024;
30'h000004ca: inst = 32'h24110080;
30'h000004cb: inst = 32'h00102021;
30'h000004cc: inst = 32'h00112821;
30'h000004cd: inst = 32'h0c0003c0;
30'h000004ce: inst = 32'h00000000;
30'h000004cf: inst = 32'h00022021;
30'h000004d0: inst = 32'h0c0001f1;
30'h000004d1: inst = 32'h00000000;
30'h000004d2: inst = 32'hafa200c0;
30'h000004d3: inst = 32'hafa200c4;
30'h000004d4: inst = 32'h8fa400c0;
30'h000004d5: inst = 32'h00000000;
30'h000004d6: inst = 32'h00102821;
30'h000004d7: inst = 32'h00113021;
30'h000004d8: inst = 32'h0c000339;
30'h000004d9: inst = 32'h00000000;
30'h000004da: inst = 32'h00022021;
30'h000004db: inst = 32'h0c000614;
30'h000004dc: inst = 32'h00000000;
30'h000004dd: inst = 32'h3c021000;
30'h000004de: inst = 32'h24441988;
30'h000004df: inst = 32'h0c000614;
30'h000004e0: inst = 32'h00000000;
30'h000004e1: inst = 32'h8fa200c4;
30'h000004e2: inst = 32'h00000000;
30'h000004e3: inst = 32'h94440000;
30'h000004e4: inst = 32'h00000000;
30'h000004e5: inst = 32'h00102821;
30'h000004e6: inst = 32'h00113021;
30'h000004e7: inst = 32'h0c0002da;
30'h000004e8: inst = 32'h00000000;
30'h000004e9: inst = 32'h080004b8;
30'h000004ea: inst = 32'h00000000;
30'h000004eb: inst = 32'h8fa400a4;
30'h000004ec: inst = 32'h00000000;
30'h000004ed: inst = 32'h3c021000;
30'h000004ee: inst = 32'h24451994;
30'h000004ef: inst = 32'h0c0005c1;
30'h000004f0: inst = 32'h00000000;
30'h000004f1: inst = 32'h14400025;
30'h000004f2: inst = 32'h00000000;
30'h000004f3: inst = 32'h3c021000;
30'h000004f4: inst = 32'h24461974;
30'h000004f5: inst = 32'h27b00024;
30'h000004f6: inst = 32'h24110080;
30'h000004f7: inst = 32'h00102021;
30'h000004f8: inst = 32'h00112821;
30'h000004f9: inst = 32'h0c0003c0;
30'h000004fa: inst = 32'h00000000;
30'h000004fb: inst = 32'h00022021;
30'h000004fc: inst = 32'h0c0001f1;
30'h000004fd: inst = 32'h00000000;
30'h000004fe: inst = 32'hafa200c8;
30'h000004ff: inst = 32'hafa200cc;
30'h00000500: inst = 32'h8fa400c8;
30'h00000501: inst = 32'h00000000;
30'h00000502: inst = 32'h00102821;
30'h00000503: inst = 32'h00113021;
30'h00000504: inst = 32'h0c000339;
30'h00000505: inst = 32'h00000000;
30'h00000506: inst = 32'h00022021;
30'h00000507: inst = 32'h0c000614;
30'h00000508: inst = 32'h00000000;
30'h00000509: inst = 32'h3c021000;
30'h0000050a: inst = 32'h24441988;
30'h0000050b: inst = 32'h0c000614;
30'h0000050c: inst = 32'h00000000;
30'h0000050d: inst = 32'h8fa200cc;
30'h0000050e: inst = 32'h00000000;
30'h0000050f: inst = 32'h90440000;
30'h00000510: inst = 32'h00000000;
30'h00000511: inst = 32'h00102821;
30'h00000512: inst = 32'h00113021;
30'h00000513: inst = 32'h0c00027b;
30'h00000514: inst = 32'h00000000;
30'h00000515: inst = 32'h080004b8;
30'h00000516: inst = 32'h00000000;
30'h00000517: inst = 32'h8fa400a4;
30'h00000518: inst = 32'h00000000;
30'h00000519: inst = 32'h3c021000;
30'h0000051a: inst = 32'h24451998;
30'h0000051b: inst = 32'h0c0005c1;
30'h0000051c: inst = 32'h00000000;
30'h0000051d: inst = 32'h1440001d;
30'h0000051e: inst = 32'h00000000;
30'h0000051f: inst = 32'h3c021000;
30'h00000520: inst = 32'h27b00024;
30'h00000521: inst = 32'h24110080;
30'h00000522: inst = 32'h24521974;
30'h00000523: inst = 32'h00102021;
30'h00000524: inst = 32'h00112821;
30'h00000525: inst = 32'h00123021;
30'h00000526: inst = 32'h0c0003c0;
30'h00000527: inst = 32'h00000000;
30'h00000528: inst = 32'h00022021;
30'h00000529: inst = 32'h0c0001f1;
30'h0000052a: inst = 32'h00000000;
30'h0000052b: inst = 32'hafa200d0;
30'h0000052c: inst = 32'h00102021;
30'h0000052d: inst = 32'h00112821;
30'h0000052e: inst = 32'h00123021;
30'h0000052f: inst = 32'h0c0003c0;
30'h00000530: inst = 32'h00000000;
30'h00000531: inst = 32'h00022021;
30'h00000532: inst = 32'h0c0001f1;
30'h00000533: inst = 32'h00000000;
30'h00000534: inst = 32'hafa200d4;
30'h00000535: inst = 32'hafa200d8;
30'h00000536: inst = 32'h8fa300d0;
30'h00000537: inst = 32'h00000000;
30'h00000538: inst = 32'hac430000;
30'h00000539: inst = 32'h08000448;
30'h0000053a: inst = 32'h00000000;
30'h0000053b: inst = 32'h8fa400a4;
30'h0000053c: inst = 32'h00000000;
30'h0000053d: inst = 32'h3c021000;
30'h0000053e: inst = 32'h2445199c;
30'h0000053f: inst = 32'h0c0005c1;
30'h00000540: inst = 32'h00000000;
30'h00000541: inst = 32'h1440001d;
30'h00000542: inst = 32'h00000000;
30'h00000543: inst = 32'h3c021000;
30'h00000544: inst = 32'h27b00024;
30'h00000545: inst = 32'h24110080;
30'h00000546: inst = 32'h24521974;
30'h00000547: inst = 32'h00102021;
30'h00000548: inst = 32'h00112821;
30'h00000549: inst = 32'h00123021;
30'h0000054a: inst = 32'h0c0003c0;
30'h0000054b: inst = 32'h00000000;
30'h0000054c: inst = 32'h00022021;
30'h0000054d: inst = 32'h0c000167;
30'h0000054e: inst = 32'h00000000;
30'h0000054f: inst = 32'ha7a200dc;
30'h00000550: inst = 32'h00102021;
30'h00000551: inst = 32'h00112821;
30'h00000552: inst = 32'h00123021;
30'h00000553: inst = 32'h0c0003c0;
30'h00000554: inst = 32'h00000000;
30'h00000555: inst = 32'h00022021;
30'h00000556: inst = 32'h0c0001f1;
30'h00000557: inst = 32'h00000000;
30'h00000558: inst = 32'hafa200e0;
30'h00000559: inst = 32'hafa200e4;
30'h0000055a: inst = 32'h97a300dc;
30'h0000055b: inst = 32'h00000000;
30'h0000055c: inst = 32'ha4430000;
30'h0000055d: inst = 32'h08000448;
30'h0000055e: inst = 32'h00000000;
30'h0000055f: inst = 32'h8fa400a4;
30'h00000560: inst = 32'h00000000;
30'h00000561: inst = 32'h3c021000;
30'h00000562: inst = 32'h244519a0;
30'h00000563: inst = 32'h0c0005c1;
30'h00000564: inst = 32'h00000000;
30'h00000565: inst = 32'h1440fee2;
30'h00000566: inst = 32'h00000000;
30'h00000567: inst = 32'h3c021000;
30'h00000568: inst = 32'h27b00024;
30'h00000569: inst = 32'h24110080;
30'h0000056a: inst = 32'h24521974;
30'h0000056b: inst = 32'h00102021;
30'h0000056c: inst = 32'h00112821;
30'h0000056d: inst = 32'h00123021;
30'h0000056e: inst = 32'h0c0003c0;
30'h0000056f: inst = 32'h00000000;
30'h00000570: inst = 32'h00022021;
30'h00000571: inst = 32'h0c0000dd;
30'h00000572: inst = 32'h00000000;
30'h00000573: inst = 32'ha3a200e8;
30'h00000574: inst = 32'h00102021;
30'h00000575: inst = 32'h00112821;
30'h00000576: inst = 32'h00123021;
30'h00000577: inst = 32'h0c0003c0;
30'h00000578: inst = 32'h00000000;
30'h00000579: inst = 32'h00022021;
30'h0000057a: inst = 32'h0c0001f1;
30'h0000057b: inst = 32'h00000000;
30'h0000057c: inst = 32'hafa200ec;
30'h0000057d: inst = 32'hafa200f0;
30'h0000057e: inst = 32'h93a300e8;
30'h0000057f: inst = 32'h00000000;
30'h00000580: inst = 32'ha0430000;
30'h00000581: inst = 32'h08000448;
30'h00000582: inst = 32'h00000000;
30'h00000583: inst = 32'h27bdffe0;
30'h00000584: inst = 32'hafa40010;
30'h00000585: inst = 32'ha3a50014;
30'h00000586: inst = 32'hafa60018;
30'h00000587: inst = 32'hafa0001c;
30'h00000588: inst = 32'h8fa2001c;
30'h00000589: inst = 32'h00000000;
30'h0000058a: inst = 32'h8fa30018;
30'h0000058b: inst = 32'h00000000;
30'h0000058c: inst = 32'h0043102b;
30'h0000058d: inst = 32'h1040000f;
30'h0000058e: inst = 32'h00000000;
30'h0000058f: inst = 32'h93a20014;
30'h00000590: inst = 32'h00000000;
30'h00000591: inst = 32'h8fa3001c;
30'h00000592: inst = 32'h00000000;
30'h00000593: inst = 32'h8fa40010;
30'h00000594: inst = 32'h00000000;
30'h00000595: inst = 32'h00831821;
30'h00000596: inst = 32'ha0620000;
30'h00000597: inst = 32'h8fa2001c;
30'h00000598: inst = 32'h00000000;
30'h00000599: inst = 32'h24420001;
30'h0000059a: inst = 32'hafa2001c;
30'h0000059b: inst = 32'h08000588;
30'h0000059c: inst = 32'h00000000;
30'h0000059d: inst = 32'h8fa20010;
30'h0000059e: inst = 32'h00000000;
30'h0000059f: inst = 32'h27bd0020;
30'h000005a0: inst = 32'h03e00008;
30'h000005a1: inst = 32'h00000000;
30'h000005a2: inst = 32'h27bdffe0;
30'h000005a3: inst = 32'hafa40010;
30'h000005a4: inst = 32'ha3a50014;
30'h000005a5: inst = 32'hafa60018;
30'h000005a6: inst = 32'hafa0001c;
30'h000005a7: inst = 32'h8fa2001c;
30'h000005a8: inst = 32'h00000000;
30'h000005a9: inst = 32'h8fa30018;
30'h000005aa: inst = 32'h00000000;
30'h000005ab: inst = 32'h0043102b;
30'h000005ac: inst = 32'h1040000f;
30'h000005ad: inst = 32'h00000000;
30'h000005ae: inst = 32'h93a20014;
30'h000005af: inst = 32'h00000000;
30'h000005b0: inst = 32'h8fa3001c;
30'h000005b1: inst = 32'h00000000;
30'h000005b2: inst = 32'h8fa40010;
30'h000005b3: inst = 32'h00000000;
30'h000005b4: inst = 32'h00831821;
30'h000005b5: inst = 32'ha0620000;
30'h000005b6: inst = 32'h8fa2001c;
30'h000005b7: inst = 32'h00000000;
30'h000005b8: inst = 32'h24420001;
30'h000005b9: inst = 32'hafa2001c;
30'h000005ba: inst = 32'h080005a7;
30'h000005bb: inst = 32'h00000000;
30'h000005bc: inst = 32'h8fa20010;
30'h000005bd: inst = 32'h00000000;
30'h000005be: inst = 32'h27bd0020;
30'h000005bf: inst = 32'h03e00008;
30'h000005c0: inst = 32'h00000000;
30'h000005c1: inst = 32'h27bdffe0;
30'h000005c2: inst = 32'hafa40014;
30'h000005c3: inst = 32'hafa50018;
30'h000005c4: inst = 32'hafa0001c;
30'h000005c5: inst = 32'h8fa20014;
30'h000005c6: inst = 32'h00000000;
30'h000005c7: inst = 32'h8fa3001c;
30'h000005c8: inst = 32'h00000000;
30'h000005c9: inst = 32'h8fa40018;
30'h000005ca: inst = 32'h00000000;
30'h000005cb: inst = 32'h00431021;
30'h000005cc: inst = 32'h00831821;
30'h000005cd: inst = 32'h80420000;
30'h000005ce: inst = 32'h00000000;
30'h000005cf: inst = 32'h80630000;
30'h000005d0: inst = 32'h00000000;
30'h000005d1: inst = 32'h10430005;
30'h000005d2: inst = 32'h00000000;
30'h000005d3: inst = 32'h24020001;
30'h000005d4: inst = 32'hafa20010;
30'h000005d5: inst = 32'h080005e7;
30'h000005d6: inst = 32'h00000000;
30'h000005d7: inst = 32'h8fa20014;
30'h000005d8: inst = 32'h00000000;
30'h000005d9: inst = 32'h8fa3001c;
30'h000005da: inst = 32'h00000000;
30'h000005db: inst = 32'h00431021;
30'h000005dc: inst = 32'h80420000;
30'h000005dd: inst = 32'h00000000;
30'h000005de: inst = 32'h10400007;
30'h000005df: inst = 32'h00000000;
30'h000005e0: inst = 32'h8fa2001c;
30'h000005e1: inst = 32'h00000000;
30'h000005e2: inst = 32'h24420001;
30'h000005e3: inst = 32'hafa2001c;
30'h000005e4: inst = 32'h080005c5;
30'h000005e5: inst = 32'h00000000;
30'h000005e6: inst = 32'hafa00010;
30'h000005e7: inst = 32'h8fa20010;
30'h000005e8: inst = 32'h00000000;
30'h000005e9: inst = 32'h27bd0020;
30'h000005ea: inst = 32'h03e00008;
30'h000005eb: inst = 32'h00000000;
30'h000005ec: inst = 32'h27bdffe8;
30'h000005ed: inst = 32'hafa40010;
30'h000005ee: inst = 32'hafa00014;
30'h000005ef: inst = 32'h8fa20010;
30'h000005f0: inst = 32'h00000000;
30'h000005f1: inst = 32'h8fa30014;
30'h000005f2: inst = 32'h00000000;
30'h000005f3: inst = 32'h00431021;
30'h000005f4: inst = 32'h80420000;
30'h000005f5: inst = 32'h00000000;
30'h000005f6: inst = 32'h10400007;
30'h000005f7: inst = 32'h00000000;
30'h000005f8: inst = 32'h8fa20014;
30'h000005f9: inst = 32'h00000000;
30'h000005fa: inst = 32'h24420001;
30'h000005fb: inst = 32'hafa20014;
30'h000005fc: inst = 32'h080005ef;
30'h000005fd: inst = 32'h00000000;
30'h000005fe: inst = 32'h8fa20014;
30'h000005ff: inst = 32'h00000000;
30'h00000600: inst = 32'h27bd0018;
30'h00000601: inst = 32'h03e00008;
30'h00000602: inst = 32'h00000000;
30'h00000603: inst = 32'h27bdffe8;
30'h00000604: inst = 32'ha3a40010;
30'h00000605: inst = 32'h3c028000;
30'h00000606: inst = 32'h34420000;
30'h00000607: inst = 32'h8c420000;
30'h00000608: inst = 32'h00000000;
30'h00000609: inst = 32'h30420001;
30'h0000060a: inst = 32'h1040fffa;
30'h0000060b: inst = 32'h00000000;
30'h0000060c: inst = 32'h3c028000;
30'h0000060d: inst = 32'h83a30010;
30'h0000060e: inst = 32'h00000000;
30'h0000060f: inst = 32'h34420008;
30'h00000610: inst = 32'hac430000;
30'h00000611: inst = 32'h27bd0018;
30'h00000612: inst = 32'h03e00008;
30'h00000613: inst = 32'h00000000;
30'h00000614: inst = 32'h27bdffd0;
30'h00000615: inst = 32'hafbf002c;
30'h00000616: inst = 32'hafa40020;
30'h00000617: inst = 32'hafa00024;
30'h00000618: inst = 32'h8fa20020;
30'h00000619: inst = 32'h00000000;
30'h0000061a: inst = 32'h8fa30024;
30'h0000061b: inst = 32'h00000000;
30'h0000061c: inst = 32'h00431021;
30'h0000061d: inst = 32'h80420000;
30'h0000061e: inst = 32'h00000000;
30'h0000061f: inst = 32'h10400010;
30'h00000620: inst = 32'h00000000;
30'h00000621: inst = 32'h8fa20020;
30'h00000622: inst = 32'h00000000;
30'h00000623: inst = 32'h8fa30024;
30'h00000624: inst = 32'h00000000;
30'h00000625: inst = 32'h00431021;
30'h00000626: inst = 32'h80440000;
30'h00000627: inst = 32'h00000000;
30'h00000628: inst = 32'h0c000603;
30'h00000629: inst = 32'h00000000;
30'h0000062a: inst = 32'h8fa20024;
30'h0000062b: inst = 32'h00000000;
30'h0000062c: inst = 32'h24420001;
30'h0000062d: inst = 32'hafa20024;
30'h0000062e: inst = 32'h08000618;
30'h0000062f: inst = 32'h00000000;
30'h00000630: inst = 32'h8fbf002c;
30'h00000631: inst = 32'h00000000;
30'h00000632: inst = 32'h27bd0030;
30'h00000633: inst = 32'h03e00008;
30'h00000634: inst = 32'h00000000;
30'h00000635: inst = 32'h27bdffd0;
30'h00000636: inst = 32'hafbf002c;
30'h00000637: inst = 32'h3c028000;
30'h00000638: inst = 32'h34420004;
30'h00000639: inst = 32'h8c420000;
30'h0000063a: inst = 32'h00000000;
30'h0000063b: inst = 32'h30420001;
30'h0000063c: inst = 32'h1040fffa;
30'h0000063d: inst = 32'h00000000;
30'h0000063e: inst = 32'h3c028000;
30'h0000063f: inst = 32'h3442000c;
30'h00000640: inst = 32'h8c420000;
30'h00000641: inst = 32'h00000000;
30'h00000642: inst = 32'ha3a20020;
30'h00000643: inst = 32'h83a20020;
30'h00000644: inst = 32'h00000000;
30'h00000645: inst = 32'h2403000d;
30'h00000646: inst = 32'h14430007;
30'h00000647: inst = 32'h00000000;
30'h00000648: inst = 32'h3c021000;
30'h00000649: inst = 32'h2444198c;
30'h0000064a: inst = 32'h0c000614;
30'h0000064b: inst = 32'h00000000;
30'h0000064c: inst = 32'h08000652;
30'h0000064d: inst = 32'h00000000;
30'h0000064e: inst = 32'h83a40020;
30'h0000064f: inst = 32'h00000000;
30'h00000650: inst = 32'h0c000603;
30'h00000651: inst = 32'h00000000;
30'h00000652: inst = 32'h83a20020;
30'h00000653: inst = 32'h00000000;
30'h00000654: inst = 32'h8fbf002c;
30'h00000655: inst = 32'h00000000;
30'h00000656: inst = 32'h27bd0030;
30'h00000657: inst = 32'h03e00008;
30'h00000658: inst = 32'h00000000;
30'h00000659: inst = 32'h0d0a0d0a;
30'h0000065a: inst = 32'h0d0a0d0a;
30'h0000065b: inst = 32'h00000000;
30'h0000065c: inst = 32'h3e200000;
30'h0000065d: inst = 32'h200d0000;
30'h0000065e: inst = 32'h66696c65;
30'h0000065f: inst = 32'h00000000;
30'h00000660: inst = 32'h6a616c00;
30'h00000661: inst = 32'h6c770000;
30'h00000662: inst = 32'h3a000000;
30'h00000663: inst = 32'h0d0a0000;
30'h00000664: inst = 32'h6c687500;
30'h00000665: inst = 32'h6c627500;
30'h00000666: inst = 32'h73770000;
30'h00000667: inst = 32'h73680000;
30'h00000668: inst = 32'h73620000;
default:      inst = 32'h00000000;
endcase
end
endmodule
