module Hazard(
  input   Clock,
  input   Reset
);

  //--|Parameters|--------------------------------------------------------------

  //--|Solution|----------------------------------------------------------------

endmodule
