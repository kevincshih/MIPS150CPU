library verilog;
use verilog.vl_types.all;
entity Datapath is
    port(
        ALUop           : in     vl_logic_vector(3 downto 0);
        REUART          : in     vl_logic;
        WEUART          : in     vl_logic;
        DinSel          : in     vl_logic;
        CTsel           : in     vl_logic;
        CTreset         : in     vl_logic;
        Stall           : in     vl_logic;
        CLK             : in     vl_logic;
        DataOutValid    : in     vl_logic;
        DataInReady     : in     vl_logic;
        reset           : in     vl_logic;
        RegWrite        : in     vl_logic;
        ICacheSel       : in     vl_logic;
        SEXTImm         : in     vl_logic;
        JRsel           : in     vl_logic;
        ControlStall    : in     vl_logic;
        PC_Sel          : in     vl_logic_vector(1 downto 0);
        ALU_Sel_A       : in     vl_logic_vector(1 downto 0);
        ALU_Sel_B       : in     vl_logic_vector(1 downto 0);
        RegDst          : in     vl_logic_vector(1 downto 0);
        UARTsel         : in     vl_logic_vector(1 downto 0);
        RDsel           : in     vl_logic_vector(1 downto 0);
        DataOut         : in     vl_logic_vector(7 downto 0);
        dcache_dout     : in     vl_logic_vector(31 downto 0);
        icache_dout     : in     vl_logic_vector(31 downto 0);
        Branch_compare  : out    vl_logic;
        RCIS            : out    vl_logic;
        offset          : out    vl_logic_vector(1 downto 0);
        Instruction     : out    vl_logic_vector(31 downto 0);
        PrevInstruction : out    vl_logic_vector(31 downto 0);
        Address         : out    vl_logic_vector(31 downto 0);
        DataOutReady    : out    vl_logic;
        DataInValid     : out    vl_logic;
        DataIn          : out    vl_logic_vector(7 downto 0);
        dcache_addr     : out    vl_logic_vector(31 downto 0);
        icache_addr     : out    vl_logic_vector(31 downto 0);
        dcache_din      : out    vl_logic_vector(31 downto 0);
        icache_din      : out    vl_logic_vector(31 downto 0);
        PC_toControl    : out    vl_logic_vector(31 downto 0);
        OldStall        : out    vl_logic
    );
end Datapath;
