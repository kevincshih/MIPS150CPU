// If #1 is in the initial block of your testbench, time advances by
// 1ns rather than 1ps
    `timescale 1ns / 1ps
    `include "Opcode.vh"
    `include "ALUop.vh"

module ControlTestbench();

parameter Halfcycle = 5; //half period is 5ns

localparam Cycle = 2 * Halfcycle;

reg Clock;

  // Clock Sinal generation:
initial Clock = 0;
always #(Halfcycle)Clock = ~Clock;

  // Register and wires
reg[31:0] Instruction;
reg[31:0] OldInstruction;
reg[31:0] Address;
reg branch;

wire RegWrite;
wire[1:0] RegDst, PCsel;
wire[1:0] AluSelA, AluSelB;
wire[3:0] ALUop, ByteSel;
wire[1:0] UARTsel, RDsel;
wire WEIM, WEDM, REUART, WEUART;

Control DUT(.Instruction(Instruction),
    .OldInstruction(OldInstruction),
	.Address(Address),
    .branch(branch),
    .reset(1'b0),
	.RegWrite(RegWrite),
    .RegDst(RegDst),
    .PCsel(PCsel),
    .AluSelA(AluSelA),
    .AluSelB(AluSelB),
    .ALUop(ALUop),
    .ByteSel(ByteSel),
    .WEIM(WEIM),
    .WEDM(WEDM),
    .REUART(REUART),
    .WEUART(WEUART),
    .UARTsel(UARTsel),
    .RDsel(RDsel));

reg[31:0] REFout;
reg[31:0] DUTout;

reg[4:0] zero = 5'b00000;
reg[4:0] s0 = 5'b10000;
reg[4:0] s1 = 5'b10001;
reg[4:0] s2 = 5'b10010;
reg[4:0] s3 = 5'b10011;
reg[15:0] imm = 16'b0;
reg[31:0] nop = 32'b0;
reg[31:0] imem = {4'b0010, 28'b0};
reg[31:0] dmem = {4'b0001, 28'b0};
reg[31:0] io = {4'b1000, 28'b0};
// Testing logic:
  
initial begin
	
	//WriteBack Logic
	$display("Write Back Logic Test");
	Instruction = {`RTYPE,s0,s0,s0,zero,`ADDU};
    OldInstruction = nop;
    Address = nop;
    branch = 1'b0;
	#1;
	if (RDsel != 2'b01) begin
	$display("FAIL: Incorrect result for RDSel expected: %h, got: %h:", 2'b01, RDsel);
	end
	if (RegDst != 2'b01) begin
	$display("FAIL: Incorrect result for RegDst expected: %h, got: %h:", 2'b01, RegDst);
	end
	#1;
	//Instruction Memory
	$display("Instruction Memory Test");
	Instruction = {`LW,s0,s0,imm};
    OldInstruction = nop;
    Address = imem;
branch = 1'b0;
	#1;
	if (WEIM != 1'b0) begin
	$display("FAIL: Incorrect result for WEIM expected: %h, got: %h:", 1'b0, WEIM);
	end
	#1;
	Instruction = {`SW,s0,s0,imm};
    OldInstruction = nop;
    Address = imem;
branch = 1'b0;
	#1;
	if (WEIM != 1'b1) begin
	$display("FAIL: Incorrect result for WEIM expected: %h, got: %h:", 1'b1, WEIM);
	end
	#1;
	
	//Data Memory
	$display("Data Memory Test");
	Instruction = {`LW,s0,s0,imm};
    OldInstruction = nop;
    Address = dmem;
branch = 1'b0;
	#1;
	if (WEDM != 1'b0) begin
	$display("FAIL: Incorrect result for WEDM expected: %h, got: %h:", 1'b0, WEDM);
	end
	if (RDsel != 2'b10) begin
	$display("FAIL: Incorrect result for RDsel expected: %h, got: %h:", 2'b10, RDsel);
	end
	#1;
	Instruction = {`SW,s0,s0,imm};
    OldInstruction = nop;
    Address = dmem;
branch = 1'b0;
	#1;
	if (WEDM != 1'b1) begin
	$display("FAIL: Incorrect result for WEDM expected: %h, got: %h:", 1'b1, WEDM);
	end
	#1;
	
	//UART I/O
	$display("UART I/O Test");
	Instruction = {`LW,s0,s0,imm};
    OldInstruction = nop;
    Address = io + 32'h0000000c;
branch = 1'b0;
	#1;
	if (REUART != 1'b1) begin
	$display("FAIL: Incorrect result for REUART expected: %h, got: %h:", 1'b1, REUART);
	end
	if (UARTsel != 2'b00) begin
	$display("FAIL: Incorrect result for UARTsel expected: %h, got: %h:", 2'b00, UARTsel);
	end
	if (RDsel != 2'b00) begin
	$display("FAIL: Incorrect result for RDsel expected: %h, got: %h:", 2'b00, RDsel);
	end	
	#1;
	
	Instruction = {`SW,s0,s0,imm};
    OldInstruction = nop;
    Address = io + 32'h8;
	#1;
	if (WEUART != 1'b1) begin
	$display("FAIL: Incorrect result for WEUART expected: %h, got: %h:", 1'b1, WEUART);
	end
	#1;
	
	//Branch/Jump Logic
	$display("Branch/Jump Test");
	Instruction = {`RTYPE,s0,zero,s0,zero,`JALR};
    	OldInstruction = nop;
    	Address = nop;
	branch = 1'b0;
	#1;
	if (PCsel != 2'b10) begin
	$display("FAIL: Incorrect result for PCSel expected: %h, got: %h:", 2'b10, PCsel);
	end
	if (AluSelA != 2'b00) begin
	$display("FAIL: Incorrect result for ALUSelA expected: %h, got: %h:", 2'b00, AluSelA);
	end
	if (AluSelB != 2'b00) begin
	$display("FAIL: Incorrect result for ALUSelB expected: %h, got: %h:", 2'b00, AluSelB);
	end
	if (RegDst != 2'b01) begin
	$display("FAIL: Incorrect result for RegDst expected: %h, got: %h:", 2'b01, RegDst);
	end
	#1;
	Instruction = {`BEQ,zero,zero,imm};
    	OldInstruction = nop;
    	Address = nop;
	branch = 1'b1;
	#1;
	if (PCsel != 2'b01) begin
	$display("FAIL: Incorrect result for PCSel expected: %h, got: %h:", 2'b01, PCsel);
	end
	if (AluSelA != 2'b01) begin
	$display("FAIL: Incorrect result for ALUSelA expected: %h, got: %h:", 2'b01, AluSelA);
	end
	if (AluSelB != 2'b01) begin
	$display("FAIL: Incorrect result for ALUSelB expected: %h, got: %h:", 2'b01, AluSelB);
	end
	#1;

	//ALU Forwarding Logic
	$display("ALU Forwarding Test");
	Instruction = {`RTYPE,s0,s0,s0,zero,`ADDU};
    	OldInstruction = {`RTYPE,s0,s0,s0,zero,`ADDU};
    	Address = nop;
	branch = 1'b0;
	#1;
	if (AluSelA != 2'b10) begin
	$display("FAIL: Incorrect result for ALUSelA expected: %h, got: %h:", 2'b10, AluSelA);
	end
	if (AluSelB != 2'b10) begin
	$display("FAIL: Incorrect result for ALUSelB expected: %h, got: %h:", 2'b10, AluSelB);
	end
	#1;
    $display("All tests passed!");
    $finish();



end
endmodule
